module leftshift1(out, shift, number);
    input shift;
    input [31:0] number;
    output [31:0] out;
    wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31;
    assign num0 = number[0];
    assign num1 = number[1];
    assign num2 = number[2];
    assign num3 = number[3];
    assign num4 = number[4];
    assign num5 = number[5];
    assign num6 = number[6];
    assign num7 = number[7];
    assign num8 = number[8];
    assign num9 = number[9];
    assign num10 = number[10];
    assign num11 = number[11];
    assign num12 = number[12];
    assign num13 = number[13];
    assign num14 = number[14];
    assign num15 = number[15];
    assign num16 = number[16];
    assign num17 = number[17];
    assign num18 = number[18];
    assign num19 = number[19];
    assign num20 = number[20];
    assign num21= number[21];
    assign num22 = number[22];
    assign num23 = number[23];
    assign num24 = number[24];
    assign num25 = number[25];
    assign num26 = number[26];
    assign num27 = number[27];
    assign num28 = number[28];
    assign num29 = number[29];
    assign num30 = number[30];
    assign num31 = number[31];

    mux_2_1 mux0(w0, shift, num0, 0);
    mux_2_1 mux1(w1, shift, num1, num0);
    mux_2_1 mux2(w2, shift, num2, num1);
    mux_2_1 mux3(w3, shift, num3, num2);
    mux_2_1 mux4(w4, shift, num4, num3);
    mux_2_1 mux5(w5, shift, num5, num4);
    mux_2_1 mux6(w6, shift, num6, num5);
    mux_2_1 mux7(w7, shift, num7, num6);
    mux_2_1 mux8(w8, shift, num8, num7);
    mux_2_1 mux9(w9, shift, num9, num8);
    mux_2_1 mux10(w10, shift, num10, num9);
    mux_2_1 mux11(w11, shift, num11, num10);
    mux_2_1 mux12(w12, shift, num12, num11);
    mux_2_1 mux13(w13, shift, num13, num12);
    mux_2_1 mux14(w14, shift, num14, num13);
    mux_2_1 mux15(w15, shift, num15, num14);
    mux_2_1 mux16(w16, shift, num16, num15);
    mux_2_1 mux17(w17, shift, num17, num16);
    mux_2_1 mux18(w18, shift, num18, num17);
    mux_2_1 mux19(w19, shift, num19, num18);
    mux_2_1 mux20(w20, shift, num20, num19);
    mux_2_1 mux21(w21, shift, num21, num20);
    mux_2_1 mux22(w22, shift, num22, num21);
    mux_2_1 mux23(w23, shift, num23, num22);
    mux_2_1 mux24(w24, shift, num24, num23);
    mux_2_1 mux25(w25, shift, num25, num24);
    mux_2_1 mux26(w26, shift, num26, num25);
    mux_2_1 mux27(w27, shift, num27, num26);
    mux_2_1 mux28(w28, shift, num28, num27);
    mux_2_1 mux29(w29, shift, num29, num28);
    mux_2_1 mux30(w30, shift, num30, num29);
    mux_2_1 mux31(w31, shift, num31, num30);

    assign out[0] = w0;
    assign out[1] = w1;
    assign out[2] = w2;
    assign out[3] = w3;
    assign out[4] = w4;
    assign out[5] = w5;
    assign out[6] = w6;
    assign out[7] = w7;
    assign out[8] = w8;
    assign out[9] = w9;
    assign out[10] = w10;
    assign out[11] = w11;
    assign out[12] = w12;
    assign out[13] = w13;
    assign out[14] = w14;
    assign out[15] = w15;
    assign out[16] = w16;
    assign out[17] = w17;
    assign out[18] = w18;
    assign out[19] = w19;
    assign out[20] = w20;
    assign out[21] = w21;
    assign out[22] = w22;
    assign out[23] = w23;
    assign out[24] = w24;
    assign out[25] = w25;
    assign out[26] = w26;
    assign out[27] = w27;
    assign out[28] = w28;
    assign out[29] = w29;
    assign out[30] = w30;
    assign out[31] = w31;
endmodule