module and32(out, A, B);
    input [31:0] A, B;
    output [31:0] out;
    
    assign num0 = A[0];
    assign num1 = A[1];
    assign num2 = A[2];
    assign num3 = A[3];
    assign num4 = A[4];
    assign num5 = A[5];
    assign num6 = A[6];
    assign num7 = A[7];
    assign num8 = A[8];
    assign num9 = A[9];
    assign num10 = A[10];
    assign num11 = A[11];
    assign num12 = A[12];
    assign num13 = A[13];
    assign num14 = A[14];
    assign num15 = A[15];
    assign num16 = A[16];
    assign num17 = A[17];
    assign num18 = A[18];
    assign num19 = A[19];
    assign num20 = A[20];
    assign num21= A[21];
    assign num22 = A[22];
    assign num23 = A[23];
    assign num24 = A[24];
    assign num25 = A[25];
    assign num26 = A[26];
    assign num27 = A[27];
    assign num28 = A[28];
    assign num29 = A[29];
    assign num30 = A[30];
    assign num31 = A[31];

    assign b0 = B[0];
    assign b1 = B[1];
    assign b2 = B[2];
    assign b3 = B[3];
    assign b4 = B[4];
    assign b5 = B[5];
    assign b6 = B[6];
    assign b7 = B[7];
    assign b8 = B[8];
    assign b9 = B[9];
    assign b10 = B[10];
    assign b11 = B[11];
    assign b12 = B[12];
    assign b13 = B[13];
    assign b14 = B[14];
    assign b15 = B[15];
    assign b16 = B[16];
    assign b17 = B[17];
    assign b18 = B[18];
    assign b19 = B[19];
    assign b20 = B[20];
    assign b21= B[21];
    assign b22 = B[22];
    assign b23 = B[23];
    assign b24 = B[24];
    assign b25 = B[25];
    assign b26 = B[26];
    assign b27 = B[27];
    assign b28 = B[28];
    assign b29 = B[29];
    assign b30 = B[30];
    assign b31 = B[31];

    wire sum0, sum1, sum2, sum3, sum4, sum5, sum6, sum7, sum8, sum9, sum10, sum11, sum12, sum13, sum14, sum15, sum16, sum17, sum18, sum19, sum20, sum21, sum22, sum23, sum24, sum25, sum26, sum27, sum28, sum29, sum30, sum31;

    and AND0(sum0, num0, b0);
    and AND1(sum1, num1, b1);
    and AND2(sum2, num2, b2);
    and AND3(sum3, num3, b3);
    and AND4(sum4, num4, b4);
    and AND5(sum5, num5, b5);
    and AND6(sum6, num6, b6);
    and AND7(sum7, num7, b7);
    and AND8(sum8, num8, b8);
    and AND9(sum9, num9, b9);
    and AND10(sum10, num10, b10);
    and AND11(sum11, num11, b11);
    and AND12(sum12, num12, b12);
    and AND13(sum13, num13, b13);
    and AND14(sum14, num14, b14);
    and AND15(sum15, num15, b15);
    and AND16(sum16, num16, b16);
    and AND17(sum17, num17, b17);
    and AND18(sum18, num18, b18);
    and AND19(sum19, num19, b19);
    and AND20(sum20, num20, b20);
    and AND21(sum21, num21, b21);
    and AND22(sum22, num22, b22);
    and AND23(sum23, num23, b23);
    and AND24(sum24, num24, b24);
    and AND25(sum25, num25, b25);
    and AND26(sum26, num26, b26);
    and AND27(sum27, num27, b27);
    and AND28(sum28, num28, b28);
    and AND29(sum29, num29, b29);
    and AND30(sum30, num30, b30);
    and AND31(sum31, num31, b31);

    assign out[0] = sum0;
    assign out[1] = sum1;
    assign out[2] = sum2;
    assign out[3] = sum3;
    assign out[4] = sum4;
    assign out[5] = sum5;
    assign out[6] = sum6;
    assign out[7] = sum7;
    assign out[8] = sum8;
    assign out[9] = sum9;
    assign out[10] = sum10;
    assign out[11] = sum11;
    assign out[12] = sum12;
    assign out[13] = sum13;
    assign out[14] = sum14;
    assign out[15] = sum15;
    assign out[16] = sum16;
    assign out[17] = sum17;
    assign out[18] = sum18;
    assign out[19] = sum19;
    assign out[20] = sum20;
    assign out[21] = sum21;
    assign out[22] = sum22;
    assign out[23] = sum23;
    assign out[24] = sum24;
    assign out[25] = sum25;
    assign out[26] = sum26;
    assign out[27] = sum27;
    assign out[28] = sum28;
    assign out[29] = sum29;
    assign out[30] = sum30;
    assign out[31] = sum31;
endmodule